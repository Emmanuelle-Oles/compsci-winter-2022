{"Models":{"obj/api/Budget.yml":[{"SourceFilePath":"obj/api/Budget.yml","FilePath":"gn231vqj.22c"}],"obj/api/Budget.Category.CategoryType.yml":[{"SourceFilePath":"obj/api/Budget.Category.CategoryType.yml","FilePath":"aakg5y2n.c1w"}],"obj/api/Budget.BudgetItemsByCategory.yml":[{"SourceFilePath":"obj/api/Budget.BudgetItemsByCategory.yml","FilePath":"o43kdvza.st4"}],"obj/api/Budget.BudgetFiles.yml":[{"SourceFilePath":"obj/api/Budget.BudgetFiles.yml","FilePath":"ui0fg0e5.3j0"}],"obj/api/Budget.BudgetItem.yml":[{"SourceFilePath":"obj/api/Budget.BudgetItem.yml","FilePath":"exytuipv.fyg"}],"obj/api/Budget.Expense.yml":[{"SourceFilePath":"obj/api/Budget.Expense.yml","FilePath":"2zqsh5fv.r2r"}],"obj/api/Budget.BudgetItemsByMonth.yml":[{"SourceFilePath":"obj/api/Budget.BudgetItemsByMonth.yml","FilePath":"a4htvyhy.oyp"}],"obj/api/Budget.Expenses.yml":[{"SourceFilePath":"obj/api/Budget.Expenses.yml","FilePath":"xth5kt02.zkd"}],"obj/api/Budget.Category.yml":[{"SourceFilePath":"obj/api/Budget.Category.yml","FilePath":"tu3bua5u.ktm"}],"obj/api/Budget.Categories.yml":[{"SourceFilePath":"obj/api/Budget.Categories.yml","FilePath":"xfofrhok.izt"}],"obj/api/Budget.HomeBudget.yml":[{"SourceFilePath":"obj/api/Budget.HomeBudget.yml","FilePath":"dg5pnukq.nyy"}]}}